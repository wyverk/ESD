-- This is the top_level VHDL file for the timer interrupt demo
-- that is being done as a hands-on demo.  The NIOS System
-- generated from the SOPC builder contains a NIOS II/s processor,
-- a 32k on-chip memory, a JTAG UART, an 8-bit output PIO that will
-- connect to the LEDs and a simple periodic interrupt 
-- generator with a 1 sec. time-out period. 

LIBRARY ieee; 
USE ieee.std_logic_1164.all; 
USE ieee.numeric_std.all;
USE ieee.std_logic_unsigned.all; 

ENTITY lab4 IS 
  port (
    

    ----- CLOCK -----
    CLOCK_50 : in std_logic;
	 
    ----- SW -----
    SW : in  std_logic_vector(9 downto 0);

    ----- KEY -----
    KEY : in std_logic_vector(3 downto 0); --for reset
	 
	 ----- LED -----
    LEDR : out  std_logic_vector(9 downto 0);  --for heartbeat
	 
	 -----?????-----
	 GPIO_0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0); --for servo pins

    ----- HEX0 ----
	 HEX0 : out std_logic_vector(6 DOWNTO 0); --for number display
	 HEX1 : out std_logic_vector(6 DOWNTO 0);
	 HEX2 : out std_logic_vector(6 DOWNTO 0);
	 HEX3 : out std_logic_vector(6 DOWNTO 0);
	 HEX4 : out std_logic_vector(6 DOWNTO 0);
	 HEX5 : out std_logic_vector(6 DOWNTO 0)
  );
  
END ENTITY;

ARCHITECTURE Structure OF lab4 IS
 
	signal reset_n : std_logic;
	signal key0_d1 : std_logic;
	signal key0_d2 : std_logic;
	signal key0_d3 : std_logic;
	
	signal key2_n : std_logic;
	signal key2_d1 : std_logic;
	signal key2_d2 : std_logic;
	signal key2_d3 : std_logic;
	
	
	signal key3_n : std_logic;
	signal key3_d1 : std_logic;
	signal key3_d2 : std_logic;
	signal key3_d3 : std_logic;
	
	signal cntr : std_logic_vector(25 downto 0);
 
	component nios_system is
		port (
			clk_clk           : in  std_logic                    := 'X';             -- clk
			reset_reset_n     : in  std_logic                    := 'X';             -- reset_n
			out_wave_out_wave : out std_logic;                                       -- out_wave
			switches_export   : in  std_logic_vector(7 downto 0) := (others => 'X'); -- export
			keys_export       : in  std_logic_vector(3 downto 0) := (others => 'X'); -- export
			hex0_export       : out std_logic_vector(6 downto 0);                    -- export
			hex1_export       : out std_logic_vector(6 downto 0);                    -- export
			hex2_export       : out std_logic_vector(6 downto 0);                    -- export
			hex3_export       : out std_logic_vector(6 downto 0);                    -- export
			hex4_export       : out std_logic_vector(6 downto 0);                    -- export
			hex5_export       : out std_logic_vector(6 downto 0)                     -- export
		);
	end component nios_system;

BEGIN 
	
	----- Syncronize the reset
  synchReset_proc : process (CLOCK_50) begin
    if (rising_edge(CLOCK_50)) then
      key0_d1 <= KEY(0);
      key0_d2 <= key0_d1;
      key0_d3 <= key0_d2;
    end if;
  end process synchReset_proc;
  reset_n <= key0_d3;
  
  
  syncKey2_proc: process(CLOCK_50)
  begin
	 if (rising_edge(CLOCK_50)) then
		key2_d1 <= KEY(2);
		key2_d2 <= key2_d1;
		key2_d3 <= key2_d2;
	 end if;
  end process;
  key2_n <= key2_d3;
  
  syncKey3_proc: process(CLOCK_50)
  begin
	 if (rising_edge(CLOCK_50)) then
		key3_d1 <= KEY(3);
		key3_d2 <= key3_d1;
		key3_d3 <= key3_d2;
	 end if;
  end process;
  key3_n <= key3_d3;
		
  --- heartbeat counter --------
  counter_proc : process (CLOCK_50) begin
    if (rising_edge(CLOCK_50)) then
      if (reset_n = '0') then
        cntr <= "00" & x"000000";
      else
        cntr <= cntr + ("00" & x"000001");
      end if;
    end if;
  end process counter_proc;
  
  LEDR(8) <= cntr(24);
	
	GPIO_0(2) <= '1';
	GPIO_0(4) <= '0';
	
-- Instantiate the Nios II system entity generated by the SOPC Builder 

	u0 : component nios_system
		port map (
			clk_clk           => CLOCK_50,           --      clk.clk
			reset_reset_n     => reset_n,     --    reset.reset_n
			out_wave_out_wave => GPIO_0(0), -- out_wave.out_wave
			switches_export   => SW(7 DOWNTO 0),   -- switches.export
			keys_export       => key3_n & key2_n & "00",       --     keys.export
			hex0_export       => HEX0,       --     hex0.export
			hex1_export       => HEX1,       --     hex1.export
			hex2_export       => HEX2,       --     hex2.export
			hex3_export       => HEX3,       --     hex3.export
			hex4_export       => HEX4,       --     hex4.export
			hex5_export       => HEX5        --     hex5.export
		);
end architecture Structure;