-- This is the top_level VHDL file for the timer interrupt demo
-- that is being done as a hands-on demo.  The NIOS System
-- generated from the SOPC builder contains a NIOS II/s processor,
-- a 32k on-chip memory, a JTAG UART, an 8-bit output PIO that will
-- connect to the LEDs and a simple periodic interrupt 
-- generator with a 1 sec. time-out period. 

LIBRARY ieee; 
USE ieee.std_logic_1164.all; 
USE ieee.numeric_std.all;
USE ieee.std_logic_unsigned.all; 

ENTITY lab3 IS 
  port (
    

    ----- CLOCK -----
    CLOCK_50 : in std_logic;
	 
    ----- SW -----
    SW : in  std_logic_vector(9 downto 0);

    ----- KEY -----
    KEY : in std_logic_vector(3 downto 0); --for reset
	 
	 ----- LED -----
    LEDR : out  std_logic_vector(9 downto 0);  --for heartbeat

    ----- HEX0 ----
	 HEX0 : out std_logic_vector(6 DOWNTO 0) --for number display
  );
  
END ENTITY;

ARCHITECTURE Structure OF lab3 IS
 
	signal reset_n : std_logic;
	signal key0_d1 : std_logic;
	signal key0_d2 : std_logic;
	signal key0_d3 : std_logic;
	signal cntr : std_logic_vector(25 downto 0);
 
	component nios_system is
		port (
			clk_clk         : in  std_logic                    := 'X';             -- clk
			reset_reset_n   : in  std_logic                    := 'X';             -- reset_n
			switches_export : in  std_logic_vector(7 downto 0) := (others => 'X'); -- export
			leds_export     : out std_logic_vector(7 downto 0);                    -- export
			hex0_export     : out std_logic_vector(6 downto 0);                    -- export
			pbs_export      : in  std_logic_vector(3 downto 0) := (others => 'X')  -- export
		);
	end component nios_system;

BEGIN 
	
	----- Syncronize the reset
  synchReset_proc : process (CLOCK_50) begin
    if (rising_edge(CLOCK_50)) then
      key0_d1 <= KEY(0);
      key0_d2 <= key0_d1;
      key0_d3 <= key0_d2;
    end if;
  end process synchReset_proc;
  reset_n <= key0_d3;
  
  --- heartbeat counter --------
  counter_proc : process (CLOCK_50) begin
    if (rising_edge(CLOCK_50)) then
      if (reset_n = '0') then
        cntr <= "00" & x"000000";
      else
        cntr <= cntr + ("00" & x"000001");
      end if;
    end if;
  end process counter_proc;
  
  LEDR(8) <= cntr(24);
	
	
-- Instantiate the Nios II system entity generated by the SOPC Builder 

	u0 : component nios_system
		port map (
			clk_clk         => CLOCK_50,         --      clk.clk
			reset_reset_n   => reset_n,   --    reset.reset_n
			switches_export => SW(7 DOWNTO 0), -- switches.export
			leds_export     => LEDR(7 DOWNTO 0),     --     leds.export
			hex0_export     => HEX0(6 DOWNTO 0),     --     hex0.export
			pbs_export      => "00" & KEY(1) & "0"  -- NIOS only has KEY1, others are dummies
		);
end architecture Structure;